`timescale 1ns / 1ps

module Counter12(
    input clk,
    output logic [3:0] q
    );
    
    always @(posedge clk) begin
        q[0] <= (!q[1] & !q[0]) | 
                ( q[1] & !q[0]) | 
                (!q[1] & !q[0]) |   
                ( q[1] & !q[0]) | 
                (!q[1] & !q[0]) | 
                ( q[1] & !q[0]); 
        
       q[1] <= (!q[1] &  q[0]) | 
               ( q[1] & !q[0]) | 
               (!q[1] &  q[0]) | 
               ( q[1] & !q[0]) | 
               (!q[1] &  q[0]) | 
               ( q[1] & !q[0]);   
       
       q[2] <= (!q[3] & !q[2] &  q[1] &  q[0]) | //0011
               (!q[3] &  q[2] & !q[1] & !q[0]) | //0100
               (!q[3] &  q[2] & !q[1] &  q[0]) | //0101
               (!q[3] &  q[2] &  q[1] & !q[0]);  //0110
       
       q[3] <= (!q[3] &  q[2] &  q[1] &  q[0]) | //0111
               ( q[3] & !q[2] & !q[1] & !q[0]) | //1000
               ( q[3] & !q[2] & !q[1] &  q[0]) | //1001
               ( q[3] & !q[2] &  q[1] & !q[0]);  //1010       
    end              
endmodule