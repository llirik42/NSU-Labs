`timescale 1ns / 1ps

module tb_fpadd();
    logic [31:0] a;
    logic [31:0] b;
    logic [31:0] s;

    fpadd DUT(.a(a), .b(b), .s(s));
    
    initial begin
        // 0 + 0
        a = 32'b00000000000000000000000000000000; b = 32'b00000000000000000000000000000000; #10; 
        
        // 0 + (-0)
        a = 32'b00000000000000000000000000000000; b = 32'b10000000000000000000000000000000; #10; 
        
        //(-0) + (-0)
        a = 32'b10000000000000000000000000000000; b = 32'b10000000000000000000000000000000; #10;
        
        // 1 + 0 
        a = 32'b00111111100000000000000000000000; b = 32'b00000000000000000000000000000000; #10; 
        
        // 1 + 1
        a = 32'b00111111100000000000000000000000; b = 32'b00111111100000000000000000000000; #10; 
        
        // 1 + (-1)
        a = 32'b00111111100000000000000000000000; b = 32'b10111111100000000000000000000000; #10; 
        
        // 1 + 0.5
        a = 32'b00111111100000000000000000000000; b = 32'b00111111000000000000000000000000; #10; 
        
        // 1 + (-0.5)
        a = 32'b00111111100000000000000000000000; b = 32'b10111111000000000000000000000000; #10; 
        
        // 0.5 + (-1)
        a = 32'b00111111000000000000000000000000; b = 32'b10111111100000000000000000000000; #10; 
        
        // 0.5 + 0.5
        a = 32'b00111111000000000000000000000000; b = 32'b00111111000000000000000000000000; #10; 
        
        // 0.5 + (-0.5)
        a = 32'b00111111000000000000000000000000; b = 32'b10111111000000000000000000000000; #10; 
        
        // 1 + 1/8
        a = 32'b00111111100000000000000000000000; b = 32'b00111110000000000000000000000000; #10; 

        // 1 - 1/8
        a = 32'b00111111100000000000000000000000; b = 32'b10111110000000000000000000000000; #10; 
     
        // (-1) + 1/8
        a = 32'b10111111100000000000000000000000; b = 32'b00111110000000000000000000000000; #10; 
     
        // 1/8 + 1/8
        a = 32'b00111110000000000000000000000000; b = 32'b00111110000000000000000000000000; #10;
     
        // 1 + 7/8
        a = 32'b00111111100000000000000000000000; b = 32'b00111111011000000000000000000000; #10; 
     
        // 1 + (-7/8)
        a = 32'b00111111100000000000000000000000; b = 32'b10111111011000000000000000000000; #10; 
        
        // 2/3 + 1/3
        a = 32'b00111110101010101010101010101011; b = 32'b00111111001010101010101010101011; #10; 
        
        // 2/3 - 1/3
        a = 32'b00111110101010101010101010101011; b = 32'b10111111001010101010101010101011; #10; 
        
        // 0.2 + 0.1
        a = 32'b00111110010011001100110011001101; b = 32'b00111101110011001100110011001101; #10; 
        
        // 0.2 - 0.1
        a = 32'b00111110010011001100110011001101; b = 32'b10111101110011001100110011001101; #10; 
        
        // 900 + 100
        a = 32'b01000100011000010000000000000000; b = 32'b01000010110010000000000000000000; #10; 
        
        // 900 - 100
        a = 32'b01000100011000010000000000000000; b = 32'b11000010110010000000000000000000; #10; 
        
        // 999 + 1
        a = 32'b01000100011110011100000000000000; b = 32'b00111111100000000000000000000000; #10; 
        
        // 999 - 1
        a = 32'b01000100011110011100000000000000; b = 32'b10111111100000000000000000000000; #10; 
 
        // max + max
        a = 32'b01111111011111111111111111111111; b = 32'b01111111011111111111111111111111; #10; 
             
        // inf + inf
        a = 32'b01111111100000000000000000000000; b = 32'b01111111100000000000000000000000; #10; 
          
        // (-inf) + (-inf)
        a = 32'b11111111100000000000000000000000; b = 32'b11111111100000000000000000000000; #10; 
          
        // inf + (-inf)
        a = 32'b01111111100000000000000000000000; b = 32'b11111111100000000000000000000000; #10; 
        
        // Nan + 0
        a = 32'b01111111110000000000000000000000; b = 32'b00000000000000000000000000000000; #10; 
        
        // Nan + 1
        a = 32'b01111111110000000000000000000000; b = 32'b00111111100000000000000000000000; #10; 
        
        // Nan + Nan
        a = 32'b01111111110000000000000000000000; b = 32'b01111111110000000000000000000000; #10; 
        
        // Nan + inf
        a = 32'b01111111110000000000000000000000; b = 32'b01111111100000000000000000000000; #10;
    $finish;
    end
endmodule
